    while odata_en = '0' loop
        idata_en <= '0';
        wait for 10 ns;
    end loop;